// jtag_axi_sys.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module jtag_axi_sys (
		output wire [7:0]  axil_master_awid,     // axil_master.awid
		output wire [31:0] axil_master_awaddr,   //            .awaddr
		output wire [7:0]  axil_master_awlen,    //            .awlen
		output wire [2:0]  axil_master_awsize,   //            .awsize
		output wire [1:0]  axil_master_awburst,  //            .awburst
		output wire [0:0]  axil_master_awlock,   //            .awlock
		output wire [3:0]  axil_master_awcache,  //            .awcache
		output wire [2:0]  axil_master_awprot,   //            .awprot
		output wire [3:0]  axil_master_awqos,    //            .awqos
		output wire [3:0]  axil_master_awregion, //            .awregion
		output wire        axil_master_awvalid,  //            .awvalid
		input  wire        axil_master_awready,  //            .awready
		output wire [31:0] axil_master_wdata,    //            .wdata
		output wire [3:0]  axil_master_wstrb,    //            .wstrb
		output wire        axil_master_wlast,    //            .wlast
		output wire        axil_master_wvalid,   //            .wvalid
		input  wire        axil_master_wready,   //            .wready
		input  wire [7:0]  axil_master_bid,      //            .bid
		input  wire [1:0]  axil_master_bresp,    //            .bresp
		input  wire        axil_master_bvalid,   //            .bvalid
		output wire        axil_master_bready,   //            .bready
		output wire [7:0]  axil_master_arid,     //            .arid
		output wire [31:0] axil_master_araddr,   //            .araddr
		output wire [7:0]  axil_master_arlen,    //            .arlen
		output wire [2:0]  axil_master_arsize,   //            .arsize
		output wire [1:0]  axil_master_arburst,  //            .arburst
		output wire [0:0]  axil_master_arlock,   //            .arlock
		output wire [3:0]  axil_master_arcache,  //            .arcache
		output wire [2:0]  axil_master_arprot,   //            .arprot
		output wire [3:0]  axil_master_arqos,    //            .arqos
		output wire [3:0]  axil_master_arregion, //            .arregion
		output wire        axil_master_arvalid,  //            .arvalid
		input  wire        axil_master_arready,  //            .arready
		input  wire [7:0]  axil_master_rid,      //            .rid
		input  wire [31:0] axil_master_rdata,    //            .rdata
		input  wire [1:0]  axil_master_rresp,    //            .rresp
		input  wire        axil_master_rlast,    //            .rlast
		input  wire        axil_master_rvalid,   //            .rvalid
		output wire        axil_master_rready,   //            .rready
		input  wire        clk_clk,              //         clk.clk
		input  wire        reset_reset_n         //       reset.reset_n
	);

	wire  [31:0] master_0_master_readdata;                   // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                    // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                       // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                 // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;              // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                      // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                  // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire   [1:0] mm_interconnect_0_axi_bridge_0_s0_awburst;  // mm_interconnect_0:axi_bridge_0_s0_awburst -> axi_bridge_0:s0_awburst
	wire   [3:0] mm_interconnect_0_axi_bridge_0_s0_arregion; // mm_interconnect_0:axi_bridge_0_s0_arregion -> axi_bridge_0:s0_arregion
	wire   [7:0] mm_interconnect_0_axi_bridge_0_s0_arlen;    // mm_interconnect_0:axi_bridge_0_s0_arlen -> axi_bridge_0:s0_arlen
	wire   [3:0] mm_interconnect_0_axi_bridge_0_s0_arqos;    // mm_interconnect_0:axi_bridge_0_s0_arqos -> axi_bridge_0:s0_arqos
	wire   [3:0] mm_interconnect_0_axi_bridge_0_s0_wstrb;    // mm_interconnect_0:axi_bridge_0_s0_wstrb -> axi_bridge_0:s0_wstrb
	wire         mm_interconnect_0_axi_bridge_0_s0_wready;   // axi_bridge_0:s0_wready -> mm_interconnect_0:axi_bridge_0_s0_wready
	wire   [7:0] mm_interconnect_0_axi_bridge_0_s0_rid;      // axi_bridge_0:s0_rid -> mm_interconnect_0:axi_bridge_0_s0_rid
	wire         mm_interconnect_0_axi_bridge_0_s0_rready;   // mm_interconnect_0:axi_bridge_0_s0_rready -> axi_bridge_0:s0_rready
	wire   [7:0] mm_interconnect_0_axi_bridge_0_s0_awlen;    // mm_interconnect_0:axi_bridge_0_s0_awlen -> axi_bridge_0:s0_awlen
	wire   [3:0] mm_interconnect_0_axi_bridge_0_s0_awqos;    // mm_interconnect_0:axi_bridge_0_s0_awqos -> axi_bridge_0:s0_awqos
	wire   [3:0] mm_interconnect_0_axi_bridge_0_s0_arcache;  // mm_interconnect_0:axi_bridge_0_s0_arcache -> axi_bridge_0:s0_arcache
	wire         mm_interconnect_0_axi_bridge_0_s0_wvalid;   // mm_interconnect_0:axi_bridge_0_s0_wvalid -> axi_bridge_0:s0_wvalid
	wire  [31:0] mm_interconnect_0_axi_bridge_0_s0_araddr;   // mm_interconnect_0:axi_bridge_0_s0_araddr -> axi_bridge_0:s0_araddr
	wire   [2:0] mm_interconnect_0_axi_bridge_0_s0_arprot;   // mm_interconnect_0:axi_bridge_0_s0_arprot -> axi_bridge_0:s0_arprot
	wire   [2:0] mm_interconnect_0_axi_bridge_0_s0_awprot;   // mm_interconnect_0:axi_bridge_0_s0_awprot -> axi_bridge_0:s0_awprot
	wire  [31:0] mm_interconnect_0_axi_bridge_0_s0_wdata;    // mm_interconnect_0:axi_bridge_0_s0_wdata -> axi_bridge_0:s0_wdata
	wire         mm_interconnect_0_axi_bridge_0_s0_arvalid;  // mm_interconnect_0:axi_bridge_0_s0_arvalid -> axi_bridge_0:s0_arvalid
	wire   [3:0] mm_interconnect_0_axi_bridge_0_s0_awcache;  // mm_interconnect_0:axi_bridge_0_s0_awcache -> axi_bridge_0:s0_awcache
	wire   [7:0] mm_interconnect_0_axi_bridge_0_s0_arid;     // mm_interconnect_0:axi_bridge_0_s0_arid -> axi_bridge_0:s0_arid
	wire   [0:0] mm_interconnect_0_axi_bridge_0_s0_arlock;   // mm_interconnect_0:axi_bridge_0_s0_arlock -> axi_bridge_0:s0_arlock
	wire   [0:0] mm_interconnect_0_axi_bridge_0_s0_awlock;   // mm_interconnect_0:axi_bridge_0_s0_awlock -> axi_bridge_0:s0_awlock
	wire  [31:0] mm_interconnect_0_axi_bridge_0_s0_awaddr;   // mm_interconnect_0:axi_bridge_0_s0_awaddr -> axi_bridge_0:s0_awaddr
	wire   [1:0] mm_interconnect_0_axi_bridge_0_s0_bresp;    // axi_bridge_0:s0_bresp -> mm_interconnect_0:axi_bridge_0_s0_bresp
	wire         mm_interconnect_0_axi_bridge_0_s0_arready;  // axi_bridge_0:s0_arready -> mm_interconnect_0:axi_bridge_0_s0_arready
	wire  [31:0] mm_interconnect_0_axi_bridge_0_s0_rdata;    // axi_bridge_0:s0_rdata -> mm_interconnect_0:axi_bridge_0_s0_rdata
	wire         mm_interconnect_0_axi_bridge_0_s0_awready;  // axi_bridge_0:s0_awready -> mm_interconnect_0:axi_bridge_0_s0_awready
	wire   [1:0] mm_interconnect_0_axi_bridge_0_s0_arburst;  // mm_interconnect_0:axi_bridge_0_s0_arburst -> axi_bridge_0:s0_arburst
	wire   [2:0] mm_interconnect_0_axi_bridge_0_s0_arsize;   // mm_interconnect_0:axi_bridge_0_s0_arsize -> axi_bridge_0:s0_arsize
	wire         mm_interconnect_0_axi_bridge_0_s0_bready;   // mm_interconnect_0:axi_bridge_0_s0_bready -> axi_bridge_0:s0_bready
	wire         mm_interconnect_0_axi_bridge_0_s0_rlast;    // axi_bridge_0:s0_rlast -> mm_interconnect_0:axi_bridge_0_s0_rlast
	wire         mm_interconnect_0_axi_bridge_0_s0_wlast;    // mm_interconnect_0:axi_bridge_0_s0_wlast -> axi_bridge_0:s0_wlast
	wire   [3:0] mm_interconnect_0_axi_bridge_0_s0_awregion; // mm_interconnect_0:axi_bridge_0_s0_awregion -> axi_bridge_0:s0_awregion
	wire   [1:0] mm_interconnect_0_axi_bridge_0_s0_rresp;    // axi_bridge_0:s0_rresp -> mm_interconnect_0:axi_bridge_0_s0_rresp
	wire   [7:0] mm_interconnect_0_axi_bridge_0_s0_awid;     // mm_interconnect_0:axi_bridge_0_s0_awid -> axi_bridge_0:s0_awid
	wire   [7:0] mm_interconnect_0_axi_bridge_0_s0_bid;      // axi_bridge_0:s0_bid -> mm_interconnect_0:axi_bridge_0_s0_bid
	wire         mm_interconnect_0_axi_bridge_0_s0_bvalid;   // axi_bridge_0:s0_bvalid -> mm_interconnect_0:axi_bridge_0_s0_bvalid
	wire   [2:0] mm_interconnect_0_axi_bridge_0_s0_awsize;   // mm_interconnect_0:axi_bridge_0_s0_awsize -> axi_bridge_0:s0_awsize
	wire         mm_interconnect_0_axi_bridge_0_s0_awvalid;  // mm_interconnect_0:axi_bridge_0_s0_awvalid -> axi_bridge_0:s0_awvalid
	wire         mm_interconnect_0_axi_bridge_0_s0_rvalid;   // axi_bridge_0:s0_rvalid -> mm_interconnect_0:axi_bridge_0_s0_rvalid
	wire         rst_controller_reset_out_reset;             // rst_controller:reset_out -> [axi_bridge_0:aresetn, mm_interconnect_0:axi_bridge_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset]

	altera_axi_bridge #(
		.USE_PIPELINE          (1),
		.USE_M0_AWID           (1),
		.USE_M0_AWREGION       (1),
		.USE_M0_AWLEN          (1),
		.USE_M0_AWSIZE         (1),
		.USE_M0_AWBURST        (1),
		.USE_M0_AWLOCK         (1),
		.USE_M0_AWCACHE        (1),
		.USE_M0_AWQOS          (1),
		.USE_S0_AWREGION       (1),
		.USE_S0_AWLOCK         (1),
		.USE_S0_AWCACHE        (1),
		.USE_S0_AWQOS          (1),
		.USE_S0_AWPROT         (1),
		.USE_M0_WSTRB          (1),
		.USE_S0_WLAST          (1),
		.USE_M0_BID            (1),
		.USE_M0_BRESP          (1),
		.USE_S0_BRESP          (1),
		.USE_M0_ARID           (1),
		.USE_M0_ARREGION       (1),
		.USE_M0_ARLEN          (1),
		.USE_M0_ARSIZE         (1),
		.USE_M0_ARBURST        (1),
		.USE_M0_ARLOCK         (1),
		.USE_M0_ARCACHE        (1),
		.USE_M0_ARQOS          (1),
		.USE_S0_ARREGION       (1),
		.USE_S0_ARLOCK         (1),
		.USE_S0_ARCACHE        (1),
		.USE_S0_ARQOS          (1),
		.USE_S0_ARPROT         (1),
		.USE_M0_RID            (1),
		.USE_M0_RRESP          (1),
		.USE_M0_RLAST          (1),
		.USE_S0_RRESP          (1),
		.M0_ID_WIDTH           (8),
		.S0_ID_WIDTH           (8),
		.DATA_WIDTH            (32),
		.WRITE_ADDR_USER_WIDTH (1),
		.READ_ADDR_USER_WIDTH  (1),
		.WRITE_DATA_USER_WIDTH (1),
		.WRITE_RESP_USER_WIDTH (1),
		.READ_DATA_USER_WIDTH  (1),
		.ADDR_WIDTH            (32),
		.USE_S0_AWUSER         (0),
		.USE_S0_ARUSER         (0),
		.USE_S0_WUSER          (0),
		.USE_S0_RUSER          (0),
		.USE_S0_BUSER          (0),
		.USE_M0_AWUSER         (0),
		.USE_M0_ARUSER         (0),
		.USE_M0_WUSER          (0),
		.USE_M0_RUSER          (0),
		.USE_M0_BUSER          (0),
		.AXI_VERSION           ("AXI4"),
		.BURST_LENGTH_WIDTH    (8),
		.LOCK_WIDTH            (1)
	) axi_bridge_0 (
		.aclk        (clk_clk),                                    //       clk.clk
		.aresetn     (~rst_controller_reset_out_reset),            // clk_reset.reset_n
		.s0_awid     (mm_interconnect_0_axi_bridge_0_s0_awid),     //        s0.awid
		.s0_awaddr   (mm_interconnect_0_axi_bridge_0_s0_awaddr),   //          .awaddr
		.s0_awlen    (mm_interconnect_0_axi_bridge_0_s0_awlen),    //          .awlen
		.s0_awsize   (mm_interconnect_0_axi_bridge_0_s0_awsize),   //          .awsize
		.s0_awburst  (mm_interconnect_0_axi_bridge_0_s0_awburst),  //          .awburst
		.s0_awlock   (mm_interconnect_0_axi_bridge_0_s0_awlock),   //          .awlock
		.s0_awcache  (mm_interconnect_0_axi_bridge_0_s0_awcache),  //          .awcache
		.s0_awprot   (mm_interconnect_0_axi_bridge_0_s0_awprot),   //          .awprot
		.s0_awqos    (mm_interconnect_0_axi_bridge_0_s0_awqos),    //          .awqos
		.s0_awregion (mm_interconnect_0_axi_bridge_0_s0_awregion), //          .awregion
		.s0_awvalid  (mm_interconnect_0_axi_bridge_0_s0_awvalid),  //          .awvalid
		.s0_awready  (mm_interconnect_0_axi_bridge_0_s0_awready),  //          .awready
		.s0_wdata    (mm_interconnect_0_axi_bridge_0_s0_wdata),    //          .wdata
		.s0_wstrb    (mm_interconnect_0_axi_bridge_0_s0_wstrb),    //          .wstrb
		.s0_wlast    (mm_interconnect_0_axi_bridge_0_s0_wlast),    //          .wlast
		.s0_wvalid   (mm_interconnect_0_axi_bridge_0_s0_wvalid),   //          .wvalid
		.s0_wready   (mm_interconnect_0_axi_bridge_0_s0_wready),   //          .wready
		.s0_bid      (mm_interconnect_0_axi_bridge_0_s0_bid),      //          .bid
		.s0_bresp    (mm_interconnect_0_axi_bridge_0_s0_bresp),    //          .bresp
		.s0_bvalid   (mm_interconnect_0_axi_bridge_0_s0_bvalid),   //          .bvalid
		.s0_bready   (mm_interconnect_0_axi_bridge_0_s0_bready),   //          .bready
		.s0_arid     (mm_interconnect_0_axi_bridge_0_s0_arid),     //          .arid
		.s0_araddr   (mm_interconnect_0_axi_bridge_0_s0_araddr),   //          .araddr
		.s0_arlen    (mm_interconnect_0_axi_bridge_0_s0_arlen),    //          .arlen
		.s0_arsize   (mm_interconnect_0_axi_bridge_0_s0_arsize),   //          .arsize
		.s0_arburst  (mm_interconnect_0_axi_bridge_0_s0_arburst),  //          .arburst
		.s0_arlock   (mm_interconnect_0_axi_bridge_0_s0_arlock),   //          .arlock
		.s0_arcache  (mm_interconnect_0_axi_bridge_0_s0_arcache),  //          .arcache
		.s0_arprot   (mm_interconnect_0_axi_bridge_0_s0_arprot),   //          .arprot
		.s0_arqos    (mm_interconnect_0_axi_bridge_0_s0_arqos),    //          .arqos
		.s0_arregion (mm_interconnect_0_axi_bridge_0_s0_arregion), //          .arregion
		.s0_arvalid  (mm_interconnect_0_axi_bridge_0_s0_arvalid),  //          .arvalid
		.s0_arready  (mm_interconnect_0_axi_bridge_0_s0_arready),  //          .arready
		.s0_rid      (mm_interconnect_0_axi_bridge_0_s0_rid),      //          .rid
		.s0_rdata    (mm_interconnect_0_axi_bridge_0_s0_rdata),    //          .rdata
		.s0_rresp    (mm_interconnect_0_axi_bridge_0_s0_rresp),    //          .rresp
		.s0_rlast    (mm_interconnect_0_axi_bridge_0_s0_rlast),    //          .rlast
		.s0_rvalid   (mm_interconnect_0_axi_bridge_0_s0_rvalid),   //          .rvalid
		.s0_rready   (mm_interconnect_0_axi_bridge_0_s0_rready),   //          .rready
		.m0_awid     (axil_master_awid),                           //        m0.awid
		.m0_awaddr   (axil_master_awaddr),                         //          .awaddr
		.m0_awlen    (axil_master_awlen),                          //          .awlen
		.m0_awsize   (axil_master_awsize),                         //          .awsize
		.m0_awburst  (axil_master_awburst),                        //          .awburst
		.m0_awlock   (axil_master_awlock),                         //          .awlock
		.m0_awcache  (axil_master_awcache),                        //          .awcache
		.m0_awprot   (axil_master_awprot),                         //          .awprot
		.m0_awqos    (axil_master_awqos),                          //          .awqos
		.m0_awregion (axil_master_awregion),                       //          .awregion
		.m0_awvalid  (axil_master_awvalid),                        //          .awvalid
		.m0_awready  (axil_master_awready),                        //          .awready
		.m0_wdata    (axil_master_wdata),                          //          .wdata
		.m0_wstrb    (axil_master_wstrb),                          //          .wstrb
		.m0_wlast    (axil_master_wlast),                          //          .wlast
		.m0_wvalid   (axil_master_wvalid),                         //          .wvalid
		.m0_wready   (axil_master_wready),                         //          .wready
		.m0_bid      (axil_master_bid),                            //          .bid
		.m0_bresp    (axil_master_bresp),                          //          .bresp
		.m0_bvalid   (axil_master_bvalid),                         //          .bvalid
		.m0_bready   (axil_master_bready),                         //          .bready
		.m0_arid     (axil_master_arid),                           //          .arid
		.m0_araddr   (axil_master_araddr),                         //          .araddr
		.m0_arlen    (axil_master_arlen),                          //          .arlen
		.m0_arsize   (axil_master_arsize),                         //          .arsize
		.m0_arburst  (axil_master_arburst),                        //          .arburst
		.m0_arlock   (axil_master_arlock),                         //          .arlock
		.m0_arcache  (axil_master_arcache),                        //          .arcache
		.m0_arprot   (axil_master_arprot),                         //          .arprot
		.m0_arqos    (axil_master_arqos),                          //          .arqos
		.m0_arregion (axil_master_arregion),                       //          .arregion
		.m0_arvalid  (axil_master_arvalid),                        //          .arvalid
		.m0_arready  (axil_master_arready),                        //          .arready
		.m0_rid      (axil_master_rid),                            //          .rid
		.m0_rdata    (axil_master_rdata),                          //          .rdata
		.m0_rresp    (axil_master_rresp),                          //          .rresp
		.m0_rlast    (axil_master_rlast),                          //          .rlast
		.m0_rvalid   (axil_master_rvalid),                         //          .rvalid
		.m0_rready   (axil_master_rready),                         //          .rready
		.s0_awuser   (1'b0),                                       // (terminated)
		.s0_wuser    (1'b0),                                       // (terminated)
		.s0_buser    (),                                           // (terminated)
		.s0_aruser   (1'b0),                                       // (terminated)
		.s0_ruser    (),                                           // (terminated)
		.m0_awuser   (),                                           // (terminated)
		.m0_wuser    (),                                           // (terminated)
		.m0_buser    (1'b0),                                       // (terminated)
		.m0_aruser   (),                                           // (terminated)
		.m0_ruser    (1'b0),                                       // (terminated)
		.m0_wid      (),                                           // (terminated)
		.s0_wid      (8'b00000000)                                 // (terminated)
	);

	jtag_axi_sys_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                       //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	jtag_axi_sys_mm_interconnect_0 mm_interconnect_0 (
		.axi_bridge_0_s0_awid                               (mm_interconnect_0_axi_bridge_0_s0_awid),     //                              axi_bridge_0_s0.awid
		.axi_bridge_0_s0_awaddr                             (mm_interconnect_0_axi_bridge_0_s0_awaddr),   //                                             .awaddr
		.axi_bridge_0_s0_awlen                              (mm_interconnect_0_axi_bridge_0_s0_awlen),    //                                             .awlen
		.axi_bridge_0_s0_awsize                             (mm_interconnect_0_axi_bridge_0_s0_awsize),   //                                             .awsize
		.axi_bridge_0_s0_awburst                            (mm_interconnect_0_axi_bridge_0_s0_awburst),  //                                             .awburst
		.axi_bridge_0_s0_awlock                             (mm_interconnect_0_axi_bridge_0_s0_awlock),   //                                             .awlock
		.axi_bridge_0_s0_awcache                            (mm_interconnect_0_axi_bridge_0_s0_awcache),  //                                             .awcache
		.axi_bridge_0_s0_awprot                             (mm_interconnect_0_axi_bridge_0_s0_awprot),   //                                             .awprot
		.axi_bridge_0_s0_awqos                              (mm_interconnect_0_axi_bridge_0_s0_awqos),    //                                             .awqos
		.axi_bridge_0_s0_awregion                           (mm_interconnect_0_axi_bridge_0_s0_awregion), //                                             .awregion
		.axi_bridge_0_s0_awvalid                            (mm_interconnect_0_axi_bridge_0_s0_awvalid),  //                                             .awvalid
		.axi_bridge_0_s0_awready                            (mm_interconnect_0_axi_bridge_0_s0_awready),  //                                             .awready
		.axi_bridge_0_s0_wdata                              (mm_interconnect_0_axi_bridge_0_s0_wdata),    //                                             .wdata
		.axi_bridge_0_s0_wstrb                              (mm_interconnect_0_axi_bridge_0_s0_wstrb),    //                                             .wstrb
		.axi_bridge_0_s0_wlast                              (mm_interconnect_0_axi_bridge_0_s0_wlast),    //                                             .wlast
		.axi_bridge_0_s0_wvalid                             (mm_interconnect_0_axi_bridge_0_s0_wvalid),   //                                             .wvalid
		.axi_bridge_0_s0_wready                             (mm_interconnect_0_axi_bridge_0_s0_wready),   //                                             .wready
		.axi_bridge_0_s0_bid                                (mm_interconnect_0_axi_bridge_0_s0_bid),      //                                             .bid
		.axi_bridge_0_s0_bresp                              (mm_interconnect_0_axi_bridge_0_s0_bresp),    //                                             .bresp
		.axi_bridge_0_s0_bvalid                             (mm_interconnect_0_axi_bridge_0_s0_bvalid),   //                                             .bvalid
		.axi_bridge_0_s0_bready                             (mm_interconnect_0_axi_bridge_0_s0_bready),   //                                             .bready
		.axi_bridge_0_s0_arid                               (mm_interconnect_0_axi_bridge_0_s0_arid),     //                                             .arid
		.axi_bridge_0_s0_araddr                             (mm_interconnect_0_axi_bridge_0_s0_araddr),   //                                             .araddr
		.axi_bridge_0_s0_arlen                              (mm_interconnect_0_axi_bridge_0_s0_arlen),    //                                             .arlen
		.axi_bridge_0_s0_arsize                             (mm_interconnect_0_axi_bridge_0_s0_arsize),   //                                             .arsize
		.axi_bridge_0_s0_arburst                            (mm_interconnect_0_axi_bridge_0_s0_arburst),  //                                             .arburst
		.axi_bridge_0_s0_arlock                             (mm_interconnect_0_axi_bridge_0_s0_arlock),   //                                             .arlock
		.axi_bridge_0_s0_arcache                            (mm_interconnect_0_axi_bridge_0_s0_arcache),  //                                             .arcache
		.axi_bridge_0_s0_arprot                             (mm_interconnect_0_axi_bridge_0_s0_arprot),   //                                             .arprot
		.axi_bridge_0_s0_arqos                              (mm_interconnect_0_axi_bridge_0_s0_arqos),    //                                             .arqos
		.axi_bridge_0_s0_arregion                           (mm_interconnect_0_axi_bridge_0_s0_arregion), //                                             .arregion
		.axi_bridge_0_s0_arvalid                            (mm_interconnect_0_axi_bridge_0_s0_arvalid),  //                                             .arvalid
		.axi_bridge_0_s0_arready                            (mm_interconnect_0_axi_bridge_0_s0_arready),  //                                             .arready
		.axi_bridge_0_s0_rid                                (mm_interconnect_0_axi_bridge_0_s0_rid),      //                                             .rid
		.axi_bridge_0_s0_rdata                              (mm_interconnect_0_axi_bridge_0_s0_rdata),    //                                             .rdata
		.axi_bridge_0_s0_rresp                              (mm_interconnect_0_axi_bridge_0_s0_rresp),    //                                             .rresp
		.axi_bridge_0_s0_rlast                              (mm_interconnect_0_axi_bridge_0_s0_rlast),    //                                             .rlast
		.axi_bridge_0_s0_rvalid                             (mm_interconnect_0_axi_bridge_0_s0_rvalid),   //                                             .rvalid
		.axi_bridge_0_s0_rready                             (mm_interconnect_0_axi_bridge_0_s0_rready),   //                                             .rready
		.clk_0_clk_clk                                      (clk_clk),                                    //                                    clk_0_clk.clk
		.axi_bridge_0_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),             // axi_bridge_0_clk_reset_reset_bridge_in_reset.reset
		.master_0_clk_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),             //     master_0_clk_reset_reset_bridge_in_reset.reset
		.master_0_master_address                            (master_0_master_address),                    //                              master_0_master.address
		.master_0_master_waitrequest                        (master_0_master_waitrequest),                //                                             .waitrequest
		.master_0_master_byteenable                         (master_0_master_byteenable),                 //                                             .byteenable
		.master_0_master_read                               (master_0_master_read),                       //                                             .read
		.master_0_master_readdata                           (master_0_master_readdata),                   //                                             .readdata
		.master_0_master_readdatavalid                      (master_0_master_readdatavalid),              //                                             .readdatavalid
		.master_0_master_write                              (master_0_master_write),                      //                                             .write
		.master_0_master_writedata                          (master_0_master_writedata)                   //                                             .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
