// aes_uart_jtag_bridge.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module aes_uart_jtag_bridge (
		input  wire  clk_clk,       //       clk.clk
		input  wire  reset_reset_n, //     reset.reset_n
		input  wire  uart_pins_rx,  // uart_pins.rx
		output wire  uart_pins_tx   //          .tx
	);

	wire  [31:0] master_0_master_readdata;                                   // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                                // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                                    // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                                       // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                                 // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                              // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                                      // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                                  // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire  [31:0] mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_awaddr;  // mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_awaddr -> aes_uart_0:s_axi_awaddr
	wire   [1:0] mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_bresp;   // aes_uart_0:s_axi_bresp -> mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_bresp
	wire         mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_arready; // aes_uart_0:s_axi_arready -> mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_arready
	wire  [31:0] mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_rdata;   // aes_uart_0:s_axi_rdata -> mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_rdata
	wire   [3:0] mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_wstrb;   // mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_wstrb -> aes_uart_0:s_axi_wstrb
	wire         mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_wready;  // aes_uart_0:s_axi_wready -> mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_wready
	wire         mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_awready; // aes_uart_0:s_axi_awready -> mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_awready
	wire         mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_rready;  // mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_rready -> aes_uart_0:s_axi_rready
	wire         mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_bready;  // mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_bready -> aes_uart_0:s_axi_bready
	wire         mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_wvalid;  // mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_wvalid -> aes_uart_0:s_axi_wvalid
	wire  [31:0] mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_araddr;  // mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_araddr -> aes_uart_0:s_axi_araddr
	wire   [2:0] mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_arprot;  // mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_arprot -> aes_uart_0:s_axi_arprot
	wire   [1:0] mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_rresp;   // aes_uart_0:s_axi_rresp -> mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_rresp
	wire   [2:0] mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_awprot;  // mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_awprot -> aes_uart_0:s_axi_awprot
	wire  [31:0] mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_wdata;   // mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_wdata -> aes_uart_0:s_axi_wdata
	wire         mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_arvalid; // mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_arvalid -> aes_uart_0:s_axi_arvalid
	wire         mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_bvalid;  // aes_uart_0:s_axi_bvalid -> mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_bvalid
	wire         mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_awvalid; // mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_awvalid -> aes_uart_0:s_axi_awvalid
	wire         mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_rvalid;  // aes_uart_0:s_axi_rvalid -> mm_interconnect_0:aes_uart_0_altera_axi4lite_slave_rvalid
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [aes_uart_0:Rst, mm_interconnect_0:aes_uart_0_reset_sink_reset_bridge_in_reset_reset]
	wire         master_0_master_reset_reset;                                // master_0:master_reset_reset -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:master_0_master_translator_reset_reset_bridge_in_reset_reset]

	AES_UART_wrapper #(
		.DATA_W (32),
		.ADDR_W (32)
	) aes_uart_0 (
		.Clk           (clk_clk),                                                    //                 clock.clk
		.s_axi_awaddr  (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_awaddr),  // altera_axi4lite_slave.awaddr
		.s_axi_awvalid (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_awvalid), //                      .awvalid
		.s_axi_awready (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_awready), //                      .awready
		.s_axi_awprot  (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_awprot),  //                      .awprot
		.s_axi_wdata   (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_wdata),   //                      .wdata
		.s_axi_wstrb   (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_wstrb),   //                      .wstrb
		.s_axi_wvalid  (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_wvalid),  //                      .wvalid
		.s_axi_wready  (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_wready),  //                      .wready
		.s_axi_bresp   (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_bresp),   //                      .bresp
		.s_axi_bvalid  (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_bvalid),  //                      .bvalid
		.s_axi_bready  (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_bready),  //                      .bready
		.s_axi_araddr  (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_araddr),  //                      .araddr
		.s_axi_arvalid (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_arvalid), //                      .arvalid
		.s_axi_arready (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_arready), //                      .arready
		.s_axi_arprot  (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_arprot),  //                      .arprot
		.s_axi_rdata   (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_rdata),   //                      .rdata
		.s_axi_rresp   (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_rresp),   //                      .rresp
		.s_axi_rvalid  (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_rvalid),  //                      .rvalid
		.s_axi_rready  (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_rready),  //                      .rready
		.Rst           (rst_controller_reset_out_reset),                             //            reset_sink.reset
		.Rx            (uart_pins_rx),                                               //           conduit_end.rx
		.Tx            (uart_pins_tx)                                                //                      .tx
	);

	aes_uart_jtag_bridge_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                       //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   (master_0_master_reset_reset)    // master_reset.reset
	);

	aes_uart_jtag_bridge_mm_interconnect_0 mm_interconnect_0 (
		.aes_uart_0_altera_axi4lite_slave_awaddr                      (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_awaddr),  //                       aes_uart_0_altera_axi4lite_slave.awaddr
		.aes_uart_0_altera_axi4lite_slave_awprot                      (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_awprot),  //                                                       .awprot
		.aes_uart_0_altera_axi4lite_slave_awvalid                     (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_awvalid), //                                                       .awvalid
		.aes_uart_0_altera_axi4lite_slave_awready                     (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_awready), //                                                       .awready
		.aes_uart_0_altera_axi4lite_slave_wdata                       (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_wdata),   //                                                       .wdata
		.aes_uart_0_altera_axi4lite_slave_wstrb                       (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_wstrb),   //                                                       .wstrb
		.aes_uart_0_altera_axi4lite_slave_wvalid                      (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_wvalid),  //                                                       .wvalid
		.aes_uart_0_altera_axi4lite_slave_wready                      (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_wready),  //                                                       .wready
		.aes_uart_0_altera_axi4lite_slave_bresp                       (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_bresp),   //                                                       .bresp
		.aes_uart_0_altera_axi4lite_slave_bvalid                      (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_bvalid),  //                                                       .bvalid
		.aes_uart_0_altera_axi4lite_slave_bready                      (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_bready),  //                                                       .bready
		.aes_uart_0_altera_axi4lite_slave_araddr                      (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_araddr),  //                                                       .araddr
		.aes_uart_0_altera_axi4lite_slave_arprot                      (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_arprot),  //                                                       .arprot
		.aes_uart_0_altera_axi4lite_slave_arvalid                     (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_arvalid), //                                                       .arvalid
		.aes_uart_0_altera_axi4lite_slave_arready                     (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_arready), //                                                       .arready
		.aes_uart_0_altera_axi4lite_slave_rdata                       (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_rdata),   //                                                       .rdata
		.aes_uart_0_altera_axi4lite_slave_rresp                       (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_rresp),   //                                                       .rresp
		.aes_uart_0_altera_axi4lite_slave_rvalid                      (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_rvalid),  //                                                       .rvalid
		.aes_uart_0_altera_axi4lite_slave_rready                      (mm_interconnect_0_aes_uart_0_altera_axi4lite_slave_rready),  //                                                       .rready
		.clk_0_clk_clk                                                (clk_clk),                                                    //                                              clk_0_clk.clk
		.aes_uart_0_reset_sink_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                             //            aes_uart_0_reset_sink_reset_bridge_in_reset.reset
		.master_0_clk_reset_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),                         //               master_0_clk_reset_reset_bridge_in_reset.reset
		.master_0_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                         // master_0_master_translator_reset_reset_bridge_in_reset.reset
		.master_0_master_address                                      (master_0_master_address),                                    //                                        master_0_master.address
		.master_0_master_waitrequest                                  (master_0_master_waitrequest),                                //                                                       .waitrequest
		.master_0_master_byteenable                                   (master_0_master_byteenable),                                 //                                                       .byteenable
		.master_0_master_read                                         (master_0_master_read),                                       //                                                       .read
		.master_0_master_readdata                                     (master_0_master_readdata),                                   //                                                       .readdata
		.master_0_master_readdatavalid                                (master_0_master_readdatavalid),                              //                                                       .readdatavalid
		.master_0_master_write                                        (master_0_master_write),                                      //                                                       .write
		.master_0_master_writedata                                    (master_0_master_writedata)                                   //                                                       .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.reset_in1      (master_0_master_reset_reset),    // reset_in1.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
